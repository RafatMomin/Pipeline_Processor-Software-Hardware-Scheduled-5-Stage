library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Pipeline_Register_N is 
   generic(N : integer := 32); 
   port( iCLK   : in std_logic;
         iRST   : in std_logic;  -- Reset signal
         i_D    : in std_logic_vector(N-1 downto 0);
         o_Q    : out std_logic_vector(N-1 downto 0));
end Pipeline_Register_N;

architecture behavioral of Pipeline_Register_N is
begin
  process(iCLK, iRST)
  begin
    if (iRST = '1') then
      o_Q <= (others => '0');  -- Reset to MIPS starting address
    elsif (rising_edge(iCLK)) then
      o_Q <= i_D;
    end if;
  end process;
end behavioral;