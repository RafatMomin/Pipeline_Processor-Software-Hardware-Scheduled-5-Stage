library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Pipeline_Register_N is 
   generic(N : integer := 32); 
   port( iCLK    : in std_logic;
         iRST    : in std_logic;  
         iSTALL  : in std_logic;  
         iFLUSH  : in std_logic;  
         i_D     : in std_logic_vector(N-1 downto 0);
         o_Q     : out std_logic_vector(N-1 downto 0));
end Pipeline_Register_N;

architecture behavioral of Pipeline_Register_N is
begin
  process(iCLK, iRST)
  begin
    if (iRST = '1') then
      o_Q <= (others => '0');  -- Reset to zeros
    elsif (rising_edge(iCLK)) then
      if (iFLUSH = '1') then
        o_Q <= (others => '0');  -- Flush/squash the register
      elsif (iSTALL = '0') then  -- Only update if not stalled
        o_Q <= i_D;
      end if;
      -- If stalled, maintain the current value
    end if;
  end process;
end behavioral;
